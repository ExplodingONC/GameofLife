// Verilog netlist created by TD v5.0.20999
// Fri Oct 16 17:59:05 2020

`timescale 1ns / 1ps
module bram_display  // bram_display.v(14)
  (
  addra,
  addrb,
  cea,
  ceb,
  clka,
  clkb,
  dia,
  dob
  );

  input [12:0] addra;  // bram_display.v(23)
  input [12:0] addrb;  // bram_display.v(24)
  input cea;  // bram_display.v(25)
  input ceb;  // bram_display.v(26)
  input clka;  // bram_display.v(27)
  input clkb;  // bram_display.v(28)
  input [23:0] dia;  // bram_display.v(22)
  output [23:0] dob;  // bram_display.v(19)

  parameter ADDR_WIDTH_A = 13;
  parameter ADDR_WIDTH_B = 13;
  parameter DATA_DEPTH_A = 8192;
  parameter DATA_DEPTH_B = 8192;
  parameter DATA_WIDTH_A = 24;
  parameter DATA_WIDTH_B = 24;
  wire [0:2] addrb_piped;
  wire  \inst_dob_mux_b0/B0_0 ;
  wire  \inst_dob_mux_b0/B0_1 ;
  wire  \inst_dob_mux_b0/B0_2 ;
  wire  \inst_dob_mux_b0/B0_3 ;
  wire  \inst_dob_mux_b0/B1_0 ;
  wire  \inst_dob_mux_b0/B1_1 ;
  wire  \inst_dob_mux_b1/B0_0 ;
  wire  \inst_dob_mux_b1/B0_1 ;
  wire  \inst_dob_mux_b1/B0_2 ;
  wire  \inst_dob_mux_b1/B0_3 ;
  wire  \inst_dob_mux_b1/B1_0 ;
  wire  \inst_dob_mux_b1/B1_1 ;
  wire  \inst_dob_mux_b10/B0_0 ;
  wire  \inst_dob_mux_b10/B0_1 ;
  wire  \inst_dob_mux_b10/B0_2 ;
  wire  \inst_dob_mux_b10/B0_3 ;
  wire  \inst_dob_mux_b10/B1_0 ;
  wire  \inst_dob_mux_b10/B1_1 ;
  wire  \inst_dob_mux_b11/B0_0 ;
  wire  \inst_dob_mux_b11/B0_1 ;
  wire  \inst_dob_mux_b11/B0_2 ;
  wire  \inst_dob_mux_b11/B0_3 ;
  wire  \inst_dob_mux_b11/B1_0 ;
  wire  \inst_dob_mux_b11/B1_1 ;
  wire  \inst_dob_mux_b12/B0_0 ;
  wire  \inst_dob_mux_b12/B0_1 ;
  wire  \inst_dob_mux_b12/B0_2 ;
  wire  \inst_dob_mux_b12/B0_3 ;
  wire  \inst_dob_mux_b12/B1_0 ;
  wire  \inst_dob_mux_b12/B1_1 ;
  wire  \inst_dob_mux_b13/B0_0 ;
  wire  \inst_dob_mux_b13/B0_1 ;
  wire  \inst_dob_mux_b13/B0_2 ;
  wire  \inst_dob_mux_b13/B0_3 ;
  wire  \inst_dob_mux_b13/B1_0 ;
  wire  \inst_dob_mux_b13/B1_1 ;
  wire  \inst_dob_mux_b14/B0_0 ;
  wire  \inst_dob_mux_b14/B0_1 ;
  wire  \inst_dob_mux_b14/B0_2 ;
  wire  \inst_dob_mux_b14/B0_3 ;
  wire  \inst_dob_mux_b14/B1_0 ;
  wire  \inst_dob_mux_b14/B1_1 ;
  wire  \inst_dob_mux_b15/B0_0 ;
  wire  \inst_dob_mux_b15/B0_1 ;
  wire  \inst_dob_mux_b15/B0_2 ;
  wire  \inst_dob_mux_b15/B0_3 ;
  wire  \inst_dob_mux_b15/B1_0 ;
  wire  \inst_dob_mux_b15/B1_1 ;
  wire  \inst_dob_mux_b16/B0_0 ;
  wire  \inst_dob_mux_b16/B0_1 ;
  wire  \inst_dob_mux_b16/B0_2 ;
  wire  \inst_dob_mux_b16/B0_3 ;
  wire  \inst_dob_mux_b16/B1_0 ;
  wire  \inst_dob_mux_b16/B1_1 ;
  wire  \inst_dob_mux_b17/B0_0 ;
  wire  \inst_dob_mux_b17/B0_1 ;
  wire  \inst_dob_mux_b17/B0_2 ;
  wire  \inst_dob_mux_b17/B0_3 ;
  wire  \inst_dob_mux_b17/B1_0 ;
  wire  \inst_dob_mux_b17/B1_1 ;
  wire  \inst_dob_mux_b2/B0_0 ;
  wire  \inst_dob_mux_b2/B0_1 ;
  wire  \inst_dob_mux_b2/B0_2 ;
  wire  \inst_dob_mux_b2/B0_3 ;
  wire  \inst_dob_mux_b2/B1_0 ;
  wire  \inst_dob_mux_b2/B1_1 ;
  wire  \inst_dob_mux_b3/B0_0 ;
  wire  \inst_dob_mux_b3/B0_1 ;
  wire  \inst_dob_mux_b3/B0_2 ;
  wire  \inst_dob_mux_b3/B0_3 ;
  wire  \inst_dob_mux_b3/B1_0 ;
  wire  \inst_dob_mux_b3/B1_1 ;
  wire  \inst_dob_mux_b4/B0_0 ;
  wire  \inst_dob_mux_b4/B0_1 ;
  wire  \inst_dob_mux_b4/B0_2 ;
  wire  \inst_dob_mux_b4/B0_3 ;
  wire  \inst_dob_mux_b4/B1_0 ;
  wire  \inst_dob_mux_b4/B1_1 ;
  wire  \inst_dob_mux_b5/B0_0 ;
  wire  \inst_dob_mux_b5/B0_1 ;
  wire  \inst_dob_mux_b5/B0_2 ;
  wire  \inst_dob_mux_b5/B0_3 ;
  wire  \inst_dob_mux_b5/B1_0 ;
  wire  \inst_dob_mux_b5/B1_1 ;
  wire  \inst_dob_mux_b6/B0_0 ;
  wire  \inst_dob_mux_b6/B0_1 ;
  wire  \inst_dob_mux_b6/B0_2 ;
  wire  \inst_dob_mux_b6/B0_3 ;
  wire  \inst_dob_mux_b6/B1_0 ;
  wire  \inst_dob_mux_b6/B1_1 ;
  wire  \inst_dob_mux_b7/B0_0 ;
  wire  \inst_dob_mux_b7/B0_1 ;
  wire  \inst_dob_mux_b7/B0_2 ;
  wire  \inst_dob_mux_b7/B0_3 ;
  wire  \inst_dob_mux_b7/B1_0 ;
  wire  \inst_dob_mux_b7/B1_1 ;
  wire  \inst_dob_mux_b8/B0_0 ;
  wire  \inst_dob_mux_b8/B0_1 ;
  wire  \inst_dob_mux_b8/B0_2 ;
  wire  \inst_dob_mux_b8/B0_3 ;
  wire  \inst_dob_mux_b8/B1_0 ;
  wire  \inst_dob_mux_b8/B1_1 ;
  wire  \inst_dob_mux_b9/B0_0 ;
  wire  \inst_dob_mux_b9/B0_1 ;
  wire  \inst_dob_mux_b9/B0_2 ;
  wire  \inst_dob_mux_b9/B0_3 ;
  wire  \inst_dob_mux_b9/B1_0 ;
  wire  \inst_dob_mux_b9/B1_1 ;
  wire inst_dob_i0_000;
  wire inst_dob_i0_001;
  wire inst_dob_i0_002;
  wire inst_dob_i0_003;
  wire inst_dob_i0_004;
  wire inst_dob_i0_005;
  wire inst_dob_i0_006;
  wire inst_dob_i0_007;
  wire inst_dob_i0_008;
  wire inst_dob_i0_009;
  wire inst_dob_i0_010;
  wire inst_dob_i0_011;
  wire inst_dob_i0_012;
  wire inst_dob_i0_013;
  wire inst_dob_i0_014;
  wire inst_dob_i0_015;
  wire inst_dob_i0_016;
  wire inst_dob_i0_017;
  wire inst_dob_i0_018;
  wire inst_dob_i0_019;
  wire inst_dob_i0_020;
  wire inst_dob_i0_021;
  wire inst_dob_i0_022;
  wire inst_dob_i0_023;
  wire inst_dob_i1_000;
  wire inst_dob_i1_001;
  wire inst_dob_i1_002;
  wire inst_dob_i1_003;
  wire inst_dob_i1_004;
  wire inst_dob_i1_005;
  wire inst_dob_i1_006;
  wire inst_dob_i1_007;
  wire inst_dob_i1_008;
  wire inst_dob_i1_009;
  wire inst_dob_i1_010;
  wire inst_dob_i1_011;
  wire inst_dob_i1_012;
  wire inst_dob_i1_013;
  wire inst_dob_i1_014;
  wire inst_dob_i1_015;
  wire inst_dob_i1_016;
  wire inst_dob_i1_017;
  wire inst_dob_i2_000;
  wire inst_dob_i2_001;
  wire inst_dob_i2_002;
  wire inst_dob_i2_003;
  wire inst_dob_i2_004;
  wire inst_dob_i2_005;
  wire inst_dob_i2_006;
  wire inst_dob_i2_007;
  wire inst_dob_i2_008;
  wire inst_dob_i2_009;
  wire inst_dob_i2_010;
  wire inst_dob_i2_011;
  wire inst_dob_i2_012;
  wire inst_dob_i2_013;
  wire inst_dob_i2_014;
  wire inst_dob_i2_015;
  wire inst_dob_i2_016;
  wire inst_dob_i2_017;
  wire inst_dob_i3_000;
  wire inst_dob_i3_001;
  wire inst_dob_i3_002;
  wire inst_dob_i3_003;
  wire inst_dob_i3_004;
  wire inst_dob_i3_005;
  wire inst_dob_i3_006;
  wire inst_dob_i3_007;
  wire inst_dob_i3_008;
  wire inst_dob_i3_009;
  wire inst_dob_i3_010;
  wire inst_dob_i3_011;
  wire inst_dob_i3_012;
  wire inst_dob_i3_013;
  wire inst_dob_i3_014;
  wire inst_dob_i3_015;
  wire inst_dob_i3_016;
  wire inst_dob_i3_017;
  wire inst_dob_i4_000;
  wire inst_dob_i4_001;
  wire inst_dob_i4_002;
  wire inst_dob_i4_003;
  wire inst_dob_i4_004;
  wire inst_dob_i4_005;
  wire inst_dob_i4_006;
  wire inst_dob_i4_007;
  wire inst_dob_i4_008;
  wire inst_dob_i4_009;
  wire inst_dob_i4_010;
  wire inst_dob_i4_011;
  wire inst_dob_i4_012;
  wire inst_dob_i4_013;
  wire inst_dob_i4_014;
  wire inst_dob_i4_015;
  wire inst_dob_i4_016;
  wire inst_dob_i4_017;
  wire inst_dob_i5_000;
  wire inst_dob_i5_001;
  wire inst_dob_i5_002;
  wire inst_dob_i5_003;
  wire inst_dob_i5_004;
  wire inst_dob_i5_005;
  wire inst_dob_i5_006;
  wire inst_dob_i5_007;
  wire inst_dob_i5_008;
  wire inst_dob_i5_009;
  wire inst_dob_i5_010;
  wire inst_dob_i5_011;
  wire inst_dob_i5_012;
  wire inst_dob_i5_013;
  wire inst_dob_i5_014;
  wire inst_dob_i5_015;
  wire inst_dob_i5_016;
  wire inst_dob_i5_017;
  wire inst_dob_i6_000;
  wire inst_dob_i6_001;
  wire inst_dob_i6_002;
  wire inst_dob_i6_003;
  wire inst_dob_i6_004;
  wire inst_dob_i6_005;
  wire inst_dob_i6_006;
  wire inst_dob_i6_007;
  wire inst_dob_i6_008;
  wire inst_dob_i6_009;
  wire inst_dob_i6_010;
  wire inst_dob_i6_011;
  wire inst_dob_i6_012;
  wire inst_dob_i6_013;
  wire inst_dob_i6_014;
  wire inst_dob_i6_015;
  wire inst_dob_i6_016;
  wire inst_dob_i6_017;
  wire inst_dob_i7_000;
  wire inst_dob_i7_001;
  wire inst_dob_i7_002;
  wire inst_dob_i7_003;
  wire inst_dob_i7_004;
  wire inst_dob_i7_005;
  wire inst_dob_i7_006;
  wire inst_dob_i7_007;
  wire inst_dob_i7_008;
  wire inst_dob_i7_009;
  wire inst_dob_i7_010;
  wire inst_dob_i7_011;
  wire inst_dob_i7_012;
  wire inst_dob_i7_013;
  wire inst_dob_i7_014;
  wire inst_dob_i7_015;
  wire inst_dob_i7_016;
  wire inst_dob_i7_017;

  assign dob[23] = inst_dob_i0_023;
  assign dob[22] = inst_dob_i0_022;
  assign dob[21] = inst_dob_i0_021;
  assign dob[20] = inst_dob_i0_020;
  assign dob[19] = inst_dob_i0_019;
  assign dob[18] = inst_dob_i0_018;
  AL_DFF_X addrb_pipe_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clkb),
    .d(addrb[10]),
    .en(ceb),
    .sr(1'b0),
    .ss(1'b0),
    .q(addrb_piped[0]));
  AL_DFF_X addrb_pipe_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clkb),
    .d(addrb[11]),
    .en(ceb),
    .sr(1'b0),
    .ss(1'b0),
    .q(addrb_piped[1]));
  AL_DFF_X addrb_pipe_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clkb),
    .d(addrb[12]),
    .en(ceb),
    .sr(1'b0),
    .ss(1'b0),
    .q(addrb_piped[2]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i0_008,inst_dob_i0_007,inst_dob_i0_006,inst_dob_i0_005,inst_dob_i0_004,inst_dob_i0_003,inst_dob_i0_002,inst_dob_i0_001,inst_dob_i0_000}));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_000000_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i0_017,inst_dob_i0_016,inst_dob_i0_015,inst_dob_i0_014,inst_dob_i0_013,inst_dob_i0_012,inst_dob_i0_011,inst_dob_i0_010,inst_dob_i0_009}));
  // address_offset=0;data_offset=18;depth=8192;width=1;num_section=1;width_per_section=1;section_size=24;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_000000_018 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n101,open_n102,open_n103,open_n104,open_n105,open_n106,open_n107,dia[18],open_n108}),
    .dob({open_n133,open_n134,open_n135,open_n136,open_n137,open_n138,open_n139,open_n140,inst_dob_i0_018}));
  // address_offset=0;data_offset=19;depth=8192;width=1;num_section=1;width_per_section=1;section_size=24;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_000000_019 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n147,open_n148,open_n149,open_n150,open_n151,open_n152,open_n153,dia[19],open_n154}),
    .dob({open_n179,open_n180,open_n181,open_n182,open_n183,open_n184,open_n185,open_n186,inst_dob_i0_019}));
  // address_offset=0;data_offset=20;depth=8192;width=1;num_section=1;width_per_section=1;section_size=24;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_000000_020 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n193,open_n194,open_n195,open_n196,open_n197,open_n198,open_n199,dia[20],open_n200}),
    .dob({open_n225,open_n226,open_n227,open_n228,open_n229,open_n230,open_n231,open_n232,inst_dob_i0_020}));
  // address_offset=0;data_offset=21;depth=8192;width=1;num_section=1;width_per_section=1;section_size=24;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_000000_021 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n239,open_n240,open_n241,open_n242,open_n243,open_n244,open_n245,dia[21],open_n246}),
    .dob({open_n271,open_n272,open_n273,open_n274,open_n275,open_n276,open_n277,open_n278,inst_dob_i0_021}));
  // address_offset=0;data_offset=22;depth=8192;width=1;num_section=1;width_per_section=1;section_size=24;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_000000_022 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n285,open_n286,open_n287,open_n288,open_n289,open_n290,open_n291,dia[22],open_n292}),
    .dob({open_n317,open_n318,open_n319,open_n320,open_n321,open_n322,open_n323,open_n324,inst_dob_i0_022}));
  // address_offset=0;data_offset=23;depth=8192;width=1;num_section=1;width_per_section=1;section_size=24;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_000000_023 (
    .addra(addra),
    .addrb(addrb),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n331,open_n332,open_n333,open_n334,open_n335,open_n336,open_n337,dia[23],open_n338}),
    .dob({open_n363,open_n364,open_n365,open_n366,open_n367,open_n368,open_n369,open_n370,inst_dob_i0_023}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i1_008,inst_dob_i1_007,inst_dob_i1_006,inst_dob_i1_005,inst_dob_i1_004,inst_dob_i1_003,inst_dob_i1_002,inst_dob_i1_001,inst_dob_i1_000}));
  // address_offset=1024;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_001024_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i1_017,inst_dob_i1_016,inst_dob_i1_015,inst_dob_i1_014,inst_dob_i1_013,inst_dob_i1_012,inst_dob_i1_011,inst_dob_i1_010,inst_dob_i1_009}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i2_008,inst_dob_i2_007,inst_dob_i2_006,inst_dob_i2_005,inst_dob_i2_004,inst_dob_i2_003,inst_dob_i2_002,inst_dob_i2_001,inst_dob_i2_000}));
  // address_offset=2048;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_002048_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i2_017,inst_dob_i2_016,inst_dob_i2_015,inst_dob_i2_014,inst_dob_i2_013,inst_dob_i2_012,inst_dob_i2_011,inst_dob_i2_010,inst_dob_i2_009}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i3_008,inst_dob_i3_007,inst_dob_i3_006,inst_dob_i3_005,inst_dob_i3_004,inst_dob_i3_003,inst_dob_i3_002,inst_dob_i3_001,inst_dob_i3_000}));
  // address_offset=3072;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_003072_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i3_017,inst_dob_i3_016,inst_dob_i3_015,inst_dob_i3_014,inst_dob_i3_013,inst_dob_i3_012,inst_dob_i3_011,inst_dob_i3_010,inst_dob_i3_009}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i4_008,inst_dob_i4_007,inst_dob_i4_006,inst_dob_i4_005,inst_dob_i4_004,inst_dob_i4_003,inst_dob_i4_002,inst_dob_i4_001,inst_dob_i4_000}));
  // address_offset=4096;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_004096_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i4_017,inst_dob_i4_016,inst_dob_i4_015,inst_dob_i4_014,inst_dob_i4_013,inst_dob_i4_012,inst_dob_i4_011,inst_dob_i4_010,inst_dob_i4_009}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i5_008,inst_dob_i5_007,inst_dob_i5_006,inst_dob_i5_005,inst_dob_i5_004,inst_dob_i5_003,inst_dob_i5_002,inst_dob_i5_001,inst_dob_i5_000}));
  // address_offset=5120;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_005120_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i5_017,inst_dob_i5_016,inst_dob_i5_015,inst_dob_i5_014,inst_dob_i5_013,inst_dob_i5_012,inst_dob_i5_011,inst_dob_i5_010,inst_dob_i5_009}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i6_008,inst_dob_i6_007,inst_dob_i6_006,inst_dob_i6_005,inst_dob_i6_004,inst_dob_i6_003,inst_dob_i6_002,inst_dob_i6_001,inst_dob_i6_000}));
  // address_offset=6144;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_006144_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i6_017,inst_dob_i6_016,inst_dob_i6_015,inst_dob_i6_014,inst_dob_i6_013,inst_dob_i6_012,inst_dob_i6_011,inst_dob_i6_010,inst_dob_i6_009}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[8:0]),
    .dob({inst_dob_i7_008,inst_dob_i7_007,inst_dob_i7_006,inst_dob_i7_005,inst_dob_i7_004,inst_dob_i7_003,inst_dob_i7_002,inst_dob_i7_001,inst_dob_i7_000}));
  // address_offset=7168;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x24_sub_007168_009 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12:10]),
    .csb(addrb[12:10]),
    .dia(dia[17:9]),
    .dob({inst_dob_i7_017,inst_dob_i7_016,inst_dob_i7_015,inst_dob_i7_014,inst_dob_i7_013,inst_dob_i7_012,inst_dob_i7_011,inst_dob_i7_010,inst_dob_i7_009}));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_0  (
    .i0(inst_dob_i0_000),
    .i1(inst_dob_i1_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_1  (
    .i0(inst_dob_i2_000),
    .i1(inst_dob_i3_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_2  (
    .i0(inst_dob_i4_000),
    .i1(inst_dob_i5_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_3  (
    .i0(inst_dob_i6_000),
    .i1(inst_dob_i7_000),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b0/B0_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b0/B0_0 ),
    .i1(\inst_dob_mux_b0/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b0/B0_2 ),
    .i1(\inst_dob_mux_b0/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b0/B1_0 ),
    .i1(\inst_dob_mux_b0/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[0]));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_0  (
    .i0(inst_dob_i0_001),
    .i1(inst_dob_i1_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_1  (
    .i0(inst_dob_i2_001),
    .i1(inst_dob_i3_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_2  (
    .i0(inst_dob_i4_001),
    .i1(inst_dob_i5_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_3  (
    .i0(inst_dob_i6_001),
    .i1(inst_dob_i7_001),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b1/B0_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b1/B0_0 ),
    .i1(\inst_dob_mux_b1/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b1/B0_2 ),
    .i1(\inst_dob_mux_b1/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b1/B1_0 ),
    .i1(\inst_dob_mux_b1/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[1]));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_0  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i1_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_1  (
    .i0(inst_dob_i2_010),
    .i1(inst_dob_i3_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_2  (
    .i0(inst_dob_i4_010),
    .i1(inst_dob_i5_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_2 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_0_3  (
    .i0(inst_dob_i6_010),
    .i1(inst_dob_i7_010),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b10/B0_3 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b10/B0_0 ),
    .i1(\inst_dob_mux_b10/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b10/B0_2 ),
    .i1(\inst_dob_mux_b10/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b10/B1_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b10/B1_0 ),
    .i1(\inst_dob_mux_b10/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[10]));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_0  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i1_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_1  (
    .i0(inst_dob_i2_011),
    .i1(inst_dob_i3_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_2  (
    .i0(inst_dob_i4_011),
    .i1(inst_dob_i5_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_2 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_0_3  (
    .i0(inst_dob_i6_011),
    .i1(inst_dob_i7_011),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b11/B0_3 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b11/B0_0 ),
    .i1(\inst_dob_mux_b11/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b11/B0_2 ),
    .i1(\inst_dob_mux_b11/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b11/B1_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b11/B1_0 ),
    .i1(\inst_dob_mux_b11/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[11]));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_0  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i1_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_1  (
    .i0(inst_dob_i2_012),
    .i1(inst_dob_i3_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_2  (
    .i0(inst_dob_i4_012),
    .i1(inst_dob_i5_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_2 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_0_3  (
    .i0(inst_dob_i6_012),
    .i1(inst_dob_i7_012),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b12/B0_3 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b12/B0_0 ),
    .i1(\inst_dob_mux_b12/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b12/B0_2 ),
    .i1(\inst_dob_mux_b12/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b12/B1_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b12/B1_0 ),
    .i1(\inst_dob_mux_b12/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[12]));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_0  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i1_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_1  (
    .i0(inst_dob_i2_013),
    .i1(inst_dob_i3_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_2  (
    .i0(inst_dob_i4_013),
    .i1(inst_dob_i5_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_2 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_0_3  (
    .i0(inst_dob_i6_013),
    .i1(inst_dob_i7_013),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b13/B0_3 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b13/B0_0 ),
    .i1(\inst_dob_mux_b13/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b13/B0_2 ),
    .i1(\inst_dob_mux_b13/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b13/B1_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b13/B1_0 ),
    .i1(\inst_dob_mux_b13/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[13]));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_0  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i1_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_1  (
    .i0(inst_dob_i2_014),
    .i1(inst_dob_i3_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_2  (
    .i0(inst_dob_i4_014),
    .i1(inst_dob_i5_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_2 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_0_3  (
    .i0(inst_dob_i6_014),
    .i1(inst_dob_i7_014),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b14/B0_3 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b14/B0_0 ),
    .i1(\inst_dob_mux_b14/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b14/B0_2 ),
    .i1(\inst_dob_mux_b14/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b14/B1_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b14/B1_0 ),
    .i1(\inst_dob_mux_b14/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[14]));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_0  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i1_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_1  (
    .i0(inst_dob_i2_015),
    .i1(inst_dob_i3_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_2  (
    .i0(inst_dob_i4_015),
    .i1(inst_dob_i5_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_2 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_0_3  (
    .i0(inst_dob_i6_015),
    .i1(inst_dob_i7_015),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b15/B0_3 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b15/B0_0 ),
    .i1(\inst_dob_mux_b15/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b15/B0_2 ),
    .i1(\inst_dob_mux_b15/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b15/B1_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b15/B1_0 ),
    .i1(\inst_dob_mux_b15/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[15]));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_0_0  (
    .i0(inst_dob_i0_016),
    .i1(inst_dob_i1_016),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b16/B0_0 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_0_1  (
    .i0(inst_dob_i2_016),
    .i1(inst_dob_i3_016),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b16/B0_1 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_0_2  (
    .i0(inst_dob_i4_016),
    .i1(inst_dob_i5_016),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b16/B0_2 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_0_3  (
    .i0(inst_dob_i6_016),
    .i1(inst_dob_i7_016),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b16/B0_3 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b16/B0_0 ),
    .i1(\inst_dob_mux_b16/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b16/B1_0 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b16/B0_2 ),
    .i1(\inst_dob_mux_b16/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b16/B1_1 ));
  AL_MUX \inst_dob_mux_b16/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b16/B1_0 ),
    .i1(\inst_dob_mux_b16/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[16]));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_0_0  (
    .i0(inst_dob_i0_017),
    .i1(inst_dob_i1_017),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b17/B0_0 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_0_1  (
    .i0(inst_dob_i2_017),
    .i1(inst_dob_i3_017),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b17/B0_1 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_0_2  (
    .i0(inst_dob_i4_017),
    .i1(inst_dob_i5_017),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b17/B0_2 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_0_3  (
    .i0(inst_dob_i6_017),
    .i1(inst_dob_i7_017),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b17/B0_3 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b17/B0_0 ),
    .i1(\inst_dob_mux_b17/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b17/B1_0 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b17/B0_2 ),
    .i1(\inst_dob_mux_b17/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b17/B1_1 ));
  AL_MUX \inst_dob_mux_b17/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b17/B1_0 ),
    .i1(\inst_dob_mux_b17/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[17]));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_0  (
    .i0(inst_dob_i0_002),
    .i1(inst_dob_i1_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_1  (
    .i0(inst_dob_i2_002),
    .i1(inst_dob_i3_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_2  (
    .i0(inst_dob_i4_002),
    .i1(inst_dob_i5_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_3  (
    .i0(inst_dob_i6_002),
    .i1(inst_dob_i7_002),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b2/B0_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b2/B0_0 ),
    .i1(\inst_dob_mux_b2/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b2/B0_2 ),
    .i1(\inst_dob_mux_b2/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b2/B1_0 ),
    .i1(\inst_dob_mux_b2/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[2]));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_0  (
    .i0(inst_dob_i0_003),
    .i1(inst_dob_i1_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_1  (
    .i0(inst_dob_i2_003),
    .i1(inst_dob_i3_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_2  (
    .i0(inst_dob_i4_003),
    .i1(inst_dob_i5_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_3  (
    .i0(inst_dob_i6_003),
    .i1(inst_dob_i7_003),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b3/B0_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b3/B0_0 ),
    .i1(\inst_dob_mux_b3/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b3/B0_2 ),
    .i1(\inst_dob_mux_b3/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b3/B1_0 ),
    .i1(\inst_dob_mux_b3/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[3]));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_0  (
    .i0(inst_dob_i0_004),
    .i1(inst_dob_i1_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_1  (
    .i0(inst_dob_i2_004),
    .i1(inst_dob_i3_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_2  (
    .i0(inst_dob_i4_004),
    .i1(inst_dob_i5_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_3  (
    .i0(inst_dob_i6_004),
    .i1(inst_dob_i7_004),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b4/B0_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b4/B0_0 ),
    .i1(\inst_dob_mux_b4/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b4/B0_2 ),
    .i1(\inst_dob_mux_b4/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b4/B1_0 ),
    .i1(\inst_dob_mux_b4/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[4]));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_0  (
    .i0(inst_dob_i0_005),
    .i1(inst_dob_i1_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_1  (
    .i0(inst_dob_i2_005),
    .i1(inst_dob_i3_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_2  (
    .i0(inst_dob_i4_005),
    .i1(inst_dob_i5_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_3  (
    .i0(inst_dob_i6_005),
    .i1(inst_dob_i7_005),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b5/B0_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b5/B0_0 ),
    .i1(\inst_dob_mux_b5/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b5/B0_2 ),
    .i1(\inst_dob_mux_b5/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b5/B1_0 ),
    .i1(\inst_dob_mux_b5/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[5]));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_0  (
    .i0(inst_dob_i0_006),
    .i1(inst_dob_i1_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_1  (
    .i0(inst_dob_i2_006),
    .i1(inst_dob_i3_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_2  (
    .i0(inst_dob_i4_006),
    .i1(inst_dob_i5_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_3  (
    .i0(inst_dob_i6_006),
    .i1(inst_dob_i7_006),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b6/B0_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b6/B0_0 ),
    .i1(\inst_dob_mux_b6/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b6/B0_2 ),
    .i1(\inst_dob_mux_b6/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b6/B1_0 ),
    .i1(\inst_dob_mux_b6/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[6]));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_0  (
    .i0(inst_dob_i0_007),
    .i1(inst_dob_i1_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_1  (
    .i0(inst_dob_i2_007),
    .i1(inst_dob_i3_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_2  (
    .i0(inst_dob_i4_007),
    .i1(inst_dob_i5_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_3  (
    .i0(inst_dob_i6_007),
    .i1(inst_dob_i7_007),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b7/B0_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b7/B0_0 ),
    .i1(\inst_dob_mux_b7/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b7/B0_2 ),
    .i1(\inst_dob_mux_b7/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b7/B1_0 ),
    .i1(\inst_dob_mux_b7/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[7]));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_0  (
    .i0(inst_dob_i0_008),
    .i1(inst_dob_i1_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_1  (
    .i0(inst_dob_i2_008),
    .i1(inst_dob_i3_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_2  (
    .i0(inst_dob_i4_008),
    .i1(inst_dob_i5_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_0_3  (
    .i0(inst_dob_i6_008),
    .i1(inst_dob_i7_008),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b8/B0_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b8/B0_0 ),
    .i1(\inst_dob_mux_b8/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b8/B0_2 ),
    .i1(\inst_dob_mux_b8/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b8/B1_0 ),
    .i1(\inst_dob_mux_b8/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[8]));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_0  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i1_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_1  (
    .i0(inst_dob_i2_009),
    .i1(inst_dob_i3_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_2  (
    .i0(inst_dob_i4_009),
    .i1(inst_dob_i5_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_2 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_0_3  (
    .i0(inst_dob_i6_009),
    .i1(inst_dob_i7_009),
    .sel(addrb_piped[0]),
    .o(\inst_dob_mux_b9/B0_3 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_dob_mux_b9/B0_0 ),
    .i1(\inst_dob_mux_b9/B0_1 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_1_1  (
    .i0(\inst_dob_mux_b9/B0_2 ),
    .i1(\inst_dob_mux_b9/B0_3 ),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b9/B1_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b9/B1_0 ),
    .i1(\inst_dob_mux_b9/B1_1 ),
    .sel(addrb_piped[2]),
    .o(dob[9]));

endmodule 

module AL_DFF_X
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_DFF u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

